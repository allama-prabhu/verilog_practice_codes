//gate level model of and gate
module AND_gt_lvl(a,b,y);
input a,b;
output y;
and(y,a,b);
endmodule


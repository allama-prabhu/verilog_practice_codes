//data flow level modeling of or gate
module ordlvl(output y, input a,b);
assign y = a | b;
endmodule


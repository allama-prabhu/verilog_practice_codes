//data flow level design for not gate
module notdlvl(output y, input a);
assign y = ~a;
endmodule


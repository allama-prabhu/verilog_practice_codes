//gate level design for not gate
module notglvl(output y, input a);
not(y,a);
endmodule


 //data flow level abstraction.
module AND_logic(y,a,b); 
input a,b;
output y;
wire y;
assign y = a & b;
endmodule


//gate level modelling of or gate
module orglvl(output y, input a,b);
or(y,a,b);
endmodule

